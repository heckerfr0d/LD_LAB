module not1(output c, input a);

nand(c, a);

endmodule

