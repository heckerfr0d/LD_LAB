module or_16(output [15:0] c, input [15:0] a, b);

or1 or_16_1 [15:0] (c, a, b);

endmodule