module and_16(output [15:0] c, input [15:0] a, b);

and1 and_16_1 [15:0] (c, a, b);

endmodule