module not_16(b, a);

output [15:0] b;
input [15:0] a;

not1 not_16_1 [15:0] (b, a);

endmodule